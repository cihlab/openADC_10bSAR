


module drc_res_2 (inout NEG, POS);

    

    PRES res_2_11 (.PRES(POS));
    PRES2 res_2_12 ();
    PRES res_2_13 (.PRES(NEG));

    PRES res_2_21 (.PRES(POS));
    PRES2 res_2_22 ();
    PRES res_2_23 (.PRES(NEG));
endmodule 



