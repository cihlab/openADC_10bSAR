
module drc_res_20 (NEG, POS);
    inout NEG;
    inout POS;
    
    PRES res_20_011 (.PRES(POS));
    PRES2 res_20_012 ();
    PRES res_20_013 (.PRES(NEG));

    PRES res_20_021 (.PRES(POS));
    PRES2 res_20_022 ();
    PRES res_20_023 (.PRES(NEG));

    PRES res_20_031 (.PRES(POS));
    PRES2 res_20_032 ();
    PRES res_20_033 (.PRES(NEG));

    PRES res_20_041 (.PRES(POS));
    PRES2 res_20_042 ();
    PRES res_20_043 (.PRES(NEG));

    PRES res_20_051 (.PRES(POS));
    PRES2 res_20_052 ();
    PRES res_20_053 (.PRES(NEG));

    PRES res_20_061 (.PRES(POS));
    PRES2 res_20_062 ();
    PRES res_20_063 (.PRES(NEG));

    PRES res_20_071 (.PRES(POS));
    PRES2 res_20_072 ();
    PRES res_20_073 (.PRES(NEG));

    PRES res_20_081 (.PRES(POS));
    PRES2 res_20_082 ();
    PRES res_20_083 (.PRES(NEG));

    PRES res_20_091 (.PRES(POS));
    PRES2 res_20_092 ();
    PRES res_20_093 (.PRES(NEG));

    PRES res_20_101 (.PRES(POS));
    PRES2 res_20_102 ();
    PRES res_20_103 (.PRES(NEG));

    PRES res_20_111 (.PRES(POS));
    PRES2 res_20_112 ();
    PRES res_20_113 (.PRES(NEG));

    PRES res_20_121 (.PRES(POS));
    PRES2 res_20_122 ();
    PRES res_20_123 (.PRES(NEG));

    PRES res_20_131 (.PRES(POS));
    PRES2 res_20_132 ();
    PRES res_20_133 (.PRES(NEG));

    PRES res_20_141 (.PRES(POS));
    PRES2 res_20_142 ();
    PRES res_20_143 (.PRES(NEG));

    PRES res_20_151 (.PRES(POS));
    PRES2 res_20_152 ();
    PRES res_20_153 (.PRES(NEG));

    PRES res_20_161 (.PRES(POS));
    PRES2 res_20_162 ();
    PRES res_20_163 (.PRES(NEG));

    PRES res_20_171 (.PRES(POS));
    PRES2 res_20_172 ();
    PRES res_20_173 (.PRES(NEG));

    PRES res_20_181 (.PRES(POS));
    PRES2 res_20_182 ();
    PRES res_20_183 (.PRES(NEG));

    PRES res_20_191 (.PRES(POS));
    PRES2 res_20_192 ();
    PRES res_20_193 (.PRES(NEG));

    PRES res_20_201 (.PRES(POS));
    PRES2 res_20_202 ();
    PRES res_20_203 (.PRES(NEG));


endmodule


