

module ADC_LP_01 (B0, B1, B10, B2, B3, B4, B5, B6, B7, B8, B9, C1, C2, C3, CLK, READY, VIN, VIP, Vdel);

    
    output B0;
    output B1;
    output B10;
    output B2;
    output B3;
    output B4;
    output B5;
    output B6;
    output B7;
    output B8;
    output B9;
    input C1;
    input C2;
    input C3;
    input CLK;
    output READY;

    input VIN;
    input VIP;



    input Vdel;

    wire net84;
    wire net117;
    wire net99;
    wire net82;
    wire net38;
    wire net37;
    wire net39;
    wire net78;
    wire net32;
    wire v8n;
    wire net50;
    wire net49;
    wire net48;
    wire net75;
    wire net45;
    wire net43;
    wire net42;
    wire v10p;
    wire net56;
    wire net55;
    wire net111;
    wire net74;
    wire net51;
    wire net95;
    wire B7p;
    wire B5p;
    wire net72;
    wire net61;
    wire net60;
    wire net59;
    wire net67;
    wire net66;
    wire net65;
    wire net64;
    wire net63;
    wire net16;
    wire net92;
    wire net77;
    wire net70;
    wire net1;
    wire net52;
    wire net58;
    wire net23;
    wire net54;
    wire net26;
    wire net68;
    wire net47;
    wire net44;
    wire net46;
    wire net57;
    wire net62;
    wire net0;
    wire net53;
    wire net102;
    wire net103;
    wire net105;
    wire net80;
    wire net107;
    wire net69;
    wire net98;
    wire c3n;
    wire net101;
    wire net100;
    wire net85;
    wire net76;
    wire net94;
    wire net93;
    wire net73;
    wire net71;
    wire net96;
    wire net79;
    wire net87;
    wire net90;
    wire c1n;
    wire net97;
    wire net89;
    wire net83;
    wire net91;
    wire net86;
    wire net81;
    wire Cal7;
    wire Cal5;
    wire Cal3;
    wire Cal6;
    wire clks;
    wire Cal4;
    wire Cal2;
    wire Cal1;
    wire Cal0;
    wire net21;
    wire net19;
    wire clk11;
    wire v2p0;
    wire v2n1;
    wire v1p0;
    wire v1n1;
    wire B1p;
    wire c2n;
    wire net88;
    wire net34;
    wire net30;
    wire net29;
    wire B4p;
    wire B3p;
    wire v9p;
    wire v7p;
    wire v5p;
    wire v2p1;
    wire v2n0;
    wire v1p1;
    wire v1n0;
    wire clkc;
    wire net113;
    wire v3p;
    wire net41;
    wire net40;
    wire net36;
    wire clk8;
    wire clk9;
    wire clk10;
    wire net17;
    wire net7;
    wire net11;
    wire outp;
    wire clk1;
    wire clk2;
    wire clk3;
    wire clk4;
    wire clk5;
    wire clk6;
    wire clk7;
    wire net4;
    wire outn;
    wire net3;
    wire B2p;
    wire net5;
    wire net6;
    wire net28;
    wire B0p;
    wire net8;
    wire net13;
    wire B9p;
    wire net14;
    wire net10;
    wire v10n;
    wire v6n;
    wire net27;
    wire v6p;
    wire B8p;
    wire net2;
    wire net12;
    wire net9;
    wire v5n;
    wire v3n;
    wire net18;
    wire net24;
    wire net20;
    wire B6p;
    wire net25;
    wire v8p;
    wire v9n;
    wire net35;
    wire net33;
    wire net15;
    wire net22;
    wire net31;
    wire v4p;
    wire v7n;
    wire v4n;

    CDAC11b_H I_18 (.CTOP(net55), .SW11(v1n1), .SW10(v1p0), .SW9(v2n1), .SW8(v2p0), .SW7(v3p), .SW6(v4p), .SW5(v5p), .SW4(v6p), .SW3(v7p), .SW2(v8p), .SW1(v9p), .SW0(v10p));
    INVD2 I_145 (.I(net88), .ZN(net85));
    DFCNQD1 I_73 (.CDN(net17), .CP(net77), .D(clk9), .Q(clk10));
    BTSW100 X0 (.CK(clks), .VIN(VIP), .VOUT(net57));
    BTSW100 X1 (.CK(clks), .VIN(VIN), .VOUT(net55));
    INVD4 I_131 (.I(net85), .ZN(B2));
    OR2D2 I_19 (.A1(outp), .A2(outn), .Z(net77));
    COMP I0 (.CALN0(Cal4), .CALN1(Cal5), .CALN2(Cal6), .CALN3(Cal7), .CALP0(Cal0), .CALP1(Cal1), .CALP2(Cal2), .CALP3(Cal3), .CLK(clkc), .OUTN(outn), .OUTP(outp), .VIN(net55), .VIP(net57));
    CDAC11b_H I_17 (.CTOP(net57), .SW11(v1n0), .SW10(v1p1), .SW9(v2n0), .SW8(v2p1), .SW7(v3n), .SW6(v4n), .SW5(v5n), .SW4(v6n), .SW3(v7n), .SW2(v8n), .SW1(v9n), .SW0(v10n));
    NR2D1 I_123 (.A1(net73), .A2(net76), .ZN(Cal5));
    DFQD1 I_92 (.CP(net86), .D(B3p), .Q(net98));
    AN3D1 I_132 (.A1(c1n), .A2(c2n), .A3(c3n), .Z(net80));
    DEL01 I_0 (.I(clk2), .Z(net3));
    INVD3 I_9 (.I(net11), .ZN(net10));
    INVD12 I_5 (.I(v2n0), .ZN(v2n1));
    INVD12 I_8 (.I(net10), .ZN(v2p0));
    AN2D1 I_2 (.A1(net3), .A2(net2), .Z(net11));
    AN2D1 I_7 (.A1(net3), .A2(B1p), .Z(net13));
    DFD1 I_1 (.CP(clk2), .D(outn), .Q(net2), .QN(B1p));
    INVD3 I_4 (.I(net13), .ZN(net4));
    INVD12 I_3 (.I(net4), .ZN(v2n0));
    INVD12 I_6 (.I(v2p0), .ZN(v2p1));
    INVD2 I_14 (.I(net12), .ZN(net7));
    AN2D1 I_27 (.A1(net15), .A2(B3p), .Z(net39));
    DEL01 I_10 (.I(clk1), .Z(net5));
    DFD1 I_11 (.CP(clk1), .D(outp), .Q(B0p), .QN(net6));
    INVD8 I_107 (.I(net70), .ZN(v4p));
    AN2D1 I_12 (.A1(net5), .A2(B0p), .Z(net12));
    AN2D1 I_13 (.A1(net5), .A2(net6), .Z(net25));
    INVD24 I_21 (.I(v1p1), .ZN(v1p0));
    DEL0 I_124 (.I(net86), .Z(net90));
    INVD24 I_15 (.I(v1n1), .ZN(v1n0));
    AN2D1 I_29 (.A1(net18), .A2(B5p), .Z(net32));
    DEL01 I_28 (.I(clk4), .Z(net15));
    INVD6 I_16 (.I(net7), .ZN(net8));
    INVD24 I_20 (.I(net8), .ZN(v1n1));
    INVD24 I_24 (.I(net9), .ZN(v1p1));
    INVD2 I_22 (.I(net25), .ZN(net31));
    DFD1 I_25 (.CP(clk4), .D(outn), .Q(net14), .QN(B3p));
    INVD6 I_23 (.I(net31), .ZN(net9));
    AN2D1 I_26 (.A1(net15), .A2(net14), .Z(net35));
    INVD2 I_106 (.I(net75), .ZN(net70));
    INVD8 I_105 (.I(net52), .ZN(v4n));
    DEL01 I_30 (.I(clk6), .Z(net18));
    AN2D1 I_31 (.A1(net18), .A2(net20), .Z(net33));
    DFD1 I_32 (.CP(clk6), .D(outn), .Q(net20), .QN(B5p));
    AN2D1 I_33 (.A1(net22), .A2(B7p), .Z(net38));
    DFD1 I_34 (.CP(clk8), .D(outn), .Q(net24), .QN(B7p));
    AN2D1 I_35 (.A1(net22), .A2(net24), .Z(net37));
    DEL01 I_36 (.I(clk8), .Z(net22));
    INVD2 I_104 (.I(net74), .ZN(net52));
    INVD4 I_103 (.I(net53), .ZN(clkc));
    DEL01 I_37 (.I(clk10), .Z(net27));
    AN2D1 I_38 (.A1(net27), .A2(net28), .Z(net43));
    DFD1 I_39 (.CP(clk10), .D(outn), .Q(net28), .QN(B9p));
    AN2D1 I_40 (.A1(net27), .A2(B9p), .Z(net42));
    INVD2 I_41 (.I(net35), .ZN(net74));
    INVD2 I_42 (.I(net39), .ZN(net75));
    INVD2 I_43 (.I(net33), .ZN(v6n));
    INVD2 I_44 (.I(net32), .ZN(v6p));
    INVD1 I_45 (.I(net38), .ZN(v8p));
    INVD1 I_46 (.I(net37), .ZN(v8n));
    INVD1 I_47 (.I(net43), .ZN(v10n));
    INVD1 I_48 (.I(net42), .ZN(v10p));
    DFD2 I_112 (.CP(net72), .D(net0), .Q(net1), .QN(net0));
    DFD1 I_49 (.CP(clk3), .D(outp), .Q(B2p), .QN(net30));
    AN2D1 I_50 (.A1(net21), .A2(B2p), .Z(net29));
    AN2D1 I_51 (.A1(net21), .A2(net30), .Z(net19));
    INVD2 I_52 (.I(net29), .ZN(net45));
    DEL01 I_53 (.I(clk3), .Z(net21));
    INVD2 I_54 (.I(net19), .ZN(net46));
    INVD4 I_55 (.I(net36), .ZN(v5n));
    DEL01 I_56 (.I(clk5), .Z(net40));
    INVD4 I_57 (.I(net34), .ZN(v5p));
    AN2D1 I_58 (.A1(net40), .A2(net41), .Z(net36));
    AN2D1 I_59 (.A1(net40), .A2(B4p), .Z(net34));
    DFD1 I_60 (.CP(clk5), .D(outp), .Q(B4p), .QN(net41));
    AN2D1 I_61 (.A1(net51), .A2(B6p), .Z(net49));
    AN2D1 I_62 (.A1(net51), .A2(net50), .Z(net48));
    INVD1 I_63 (.I(net49), .ZN(v7p));
    DEL01 I_64 (.I(clk7), .Z(net51));
    DFD1 I_65 (.CP(clk7), .D(outp), .Q(B6p), .QN(net50));
    INVD1 I_66 (.I(net48), .ZN(v7n));
    INVD1 I_67 (.I(net59), .ZN(v9n));
    DFD1 I_68 (.CP(clk9), .D(outp), .Q(B8p), .QN(net56));
    TIEH I_101 (.Z(net44));
    DEL01 I_69 (.I(clk9), .Z(net61));
    INVD1 I_70 (.I(net60), .ZN(v9p));
    AN2D1 I_71 (.A1(net61), .A2(net56), .Z(net59));
    AN2D1 I_72 (.A1(net61), .A2(B8p), .Z(net60));
    DFCNQD1 I_74 (.CDN(net17), .CP(net77), .D(clk8), .Q(clk9));
    DFCNQD1 I_75 (.CDN(net17), .CP(net77), .D(clk7), .Q(clk8));
    DFCNQD1 I_76 (.CDN(net17), .CP(net77), .D(clk6), .Q(clk7));
    DFCNQD1 I_77 (.CDN(net17), .CP(net77), .D(clk5), .Q(clk6));
    DFCNQD1 I_78 (.CDN(net17), .CP(net77), .D(net44), .Q(clk1));
    INVD4 I_79 (.I(clks), .ZN(net17));
    INVD1 I_87 (.I(net63), .ZN(net16));
    VCDC2 X2 (.CK(net16), .TL(net66), .VIN(Vdel), .ZN(net65));
    VCDC2 X3 (.CK(net77), .TL(net64), .VIN(Vdel), .ZN(net63));
    DFQD1 I_94 (.CP(net86), .D(B2p), .Q(net99));
    DFQD1 I_95 (.CP(net86), .D(B5p), .Q(net95));
    DFQD1 I_96 (.CP(net86), .D(B6p), .Q(net91));
    DFQD1 I_97 (.CP(net86), .D(B7p), .Q(net89));
    DFCNQD1 I_80 (.CDN(net17), .CP(net77), .D(clk4), .Q(clk5));
    DFCNQD1 I_81 (.CDN(net17), .CP(net77), .D(clk3), .Q(clk4));
    DFCNQD1 I_82 (.CDN(net17), .CP(net77), .D(clk2), .Q(clk3));
    DFCNQD1 I_83 (.CDN(net17), .CP(net77), .D(clk1), .Q(clk2));
    DFQD1 I_91 (.CP(net86), .D(B1p), .Q(net101));
    NR2D1 I_122 (.A1(net81), .A2(net82), .ZN(Cal3));
    DFQD1 I_93 (.CP(net86), .D(B4p), .Q(net97));
    INVD1 I_102 (.I(net58), .ZN(net53));
    DFQD1 I_90 (.CP(net86), .D(B0p), .Q(net103));
    INVD2 I_88 (.I(clk11), .ZN(net26));
    INVD4 I_89 (.I(net26), .ZN(net86));
    INVD1 I_86 (.I(net65), .ZN(net67));
    DFCNQD1 I_84 (.CDN(net17), .CP(net77), .D(clk10), .Q(clk11));
    NR3D0 I_85 (.A1(clk11), .A2(net67), .A3(clks), .ZN(net58));
    DFQD1 I_98 (.CP(net86), .D(B8p), .Q(net88));
    DFQD1 I_99 (.CP(net86), .D(B9p), .Q(net84));
    INVD4 I_108 (.I(net45), .ZN(net62));
    CKBD3 I_115 (.I(CLK), .Z(net72));
    AN2D2 I_114 (.A1(net1), .A2(net54), .Z(clks));
    INVD8 I_109 (.I(net62), .ZN(v3p));
    INVD4 I_110 (.I(net46), .ZN(net78));
    INVD8 I_111 (.I(net78), .ZN(v3n));
    DEL4 I_113 (.I(net72), .Z(net54));
    DFQD1 I_100 (.CP(net86), .D(outp), .Q(net23));
    INVD1 I_120 (.I(C2), .ZN(c2n));
    INVD1 I_121 (.I(C3), .ZN(c3n));
    INVD1 I_119 (.I(C1), .ZN(c1n));
    ND3D1 I_118 (.A1(C1), .A2(C2), .A3(C3), .ZN(Cal1));
    ND2D1 I_117 (.A1(C1), .A2(C2), .ZN(Cal2));
    AN2D1 I_116 (.A1(C2), .A2(C1), .Z(net81));
    INVD4 I_130 (.I(net83), .ZN(B0));
    INVD2 I_129 (.I(net23), .ZN(net83));
    AN3D1 I_133 (.A1(C1), .A2(c2n), .A3(c3n), .Z(net73));
    AN3D1 I_134 (.A1(c1n), .A2(C2), .A3(C3), .Z(net76));
    OR3D1 I_135 (.A1(net80), .A2(net79), .A3(net71), .Z(Cal7));
    OR3D1 I_136 (.A1(net68), .A2(net69), .A3(net47), .Z(Cal6));
    AN2D1 I_137 (.A1(C1), .A2(C3), .Z(net82));
    AN2D1 I_138 (.A1(C2), .A2(C1), .Z(net79));
    AN2D1 I_139 (.A1(C1), .A2(C3), .Z(net71));
    AN2D1 I_140 (.A1(c1n), .A2(c2n), .Z(net68));
    AN2D1 I_141 (.A1(C2), .A2(C1), .Z(net69));
    AN2D1 I_142 (.A1(C1), .A2(C3), .Z(net47));
    ND3D1 I_143 (.A1(C1), .A2(c2n), .A3(c3n), .ZN(Cal4));
    INVD8 I_128 (.I(net92), .ZN(READY));
    INVD3 I_127 (.I(net87), .ZN(net92));
    DEL0 I_126 (.I(net94), .Z(net87));
    DEL0 I_125 (.I(net90), .Z(net94));
    TIEH I_144 (.Z(Cal0));
    INVD2 I_146 (.I(net91), .ZN(net93));
    INVD4 I_147 (.I(net93), .ZN(B4));
    INVD4 I_148 (.I(net96), .ZN(B6));
    INVD2 I_149 (.I(net97), .ZN(net96));
    INVD2 I_150 (.I(net99), .ZN(net100));
    INVD4 I_151 (.I(net100), .ZN(B8));
    INVD4 I_152 (.I(net102), .ZN(B10));
    INVD2 I_153 (.I(net103), .ZN(net102));
    INVD4 I_154 (.I(net107), .ZN(B3));
    INVD4 I_155 (.I(net105), .ZN(B5));
    INVD2 I_156 (.I(net89), .ZN(net107));
    INVD2 I_157 (.I(net95), .ZN(net105));
    INVD4 I_158 (.I(net113), .ZN(B7));
    INVD4 I_159 (.I(net111), .ZN(B9));
    INVD2 I_160 (.I(net98), .ZN(net113));
    INVD2 I_161 (.I(net101), .ZN(net111));
    INVD2 I_164 (.I(net84), .ZN(net117));
    INVD4 I_165 (.I(net117), .ZN(B1));
endmodule // ADC_LP_01_netlist


